`include "tb_drv_common.sv"
`include "tb_drv_axi.sv"
`include "tb_drv_axis.sv"