`ifndef TB_DEF_SV
`define TB_DEF_SV

`endif
